parameter WR_PTR_WIDTH = 4;
parameter RD_PTR_WIDTH = 4;
parameter ADDR_WIDTH = 4;
parameter DATA_WIDTH = 4;
